library verilog;
use verilog.vl_types.all;
entity Testef2_vlg_vec_tst is
end Testef2_vlg_vec_tst;
