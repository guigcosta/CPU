library verilog;
use verilog.vl_types.all;
entity Teste2_vlg_vec_tst is
end Teste2_vlg_vec_tst;
